module notgate(
    input a,
    output b
);

// Assign the NOT operation to output b
assign b = ~a;

endmodule
